
module Lego_control_unit #()(

);

endmodule