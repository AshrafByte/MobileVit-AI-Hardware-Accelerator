//==============================================================================
// Package: accelerator_pkg
// Description: Main package for MobileVit AI Hardware Accelerator
//              Imports all sub-packages for convenience
// Author: MobileVit Team
// Date: October 9, 2025
//==============================================================================

package accelerator_pkg;

    // Import all sub-packages
    import accelerator_common_pkg::*;
    import accelerator_matmul_pkg::*;
    import accelerator_norm_pkg::*;
    import accelerator_activation_pkg::*;

endpackage : accelerator_pkg
